** sch_path: /home/jrsharp/home_mnt/asic/iic-jku-analog/2_1_1-Large-signal-MOSFET-Model/nmos-sweep.sch
**.subckt nmos-sweep


* model can be e.g. sky130_fd_pr__nfet_01v8 
XM1 net_ds net_gs GND GND ${MODEL} L=${LENGTH} W=${WIDTH} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vds net1 GND 1.8
Vd net1 net_ds 0
.save i(vd)
Vgs net_gs GND 0.8
**** begin user architecture code

.lib /home/jrsharp/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt


.temp 27
.control
save all
save @m.XM1.m${MODEL}[id]
save @m.XM1.m${MODEL}[gm]
save @m.XM1.m${MODEL}[gds]
save @m.XM1.m${MODEL}[vth]
save @m.XM1.m${MODEL}[cgg]
save @m.XM1.m${MODEL}[cgd]
save @m.XM1.m${MODEL}[vdss]
save @m.XM1.m${MODEL}[fug]
save @m.XM1.m${MODEL}[rg]
save @m.XM1.m${MODEL}[sid]
op
write ${FILE}
set appendwrite
dc Vds 0 1.8 0.01 Vgs 0 1.8 0.1
write ${FILE}
quit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
